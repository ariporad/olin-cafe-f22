`ifndef INITIAL_CONDITIONS
`define INITIAL_CONDITIONS

`define INIT_5x5_PERIOD2_TOAD { \
  7'b0000000, \
  7'b0010000, \
  7'b0011000, \
  7'b0011000, \
  7'b0001000, \
  7'b0000000, \
  7'b0000000 \
}

`define INIT_5x5_PERIOD2_BLINKER { \
  7'b0000000, \
  7'b0000000, \
  7'b0000000, \
  7'b0011100, \
  7'b0000000, \
  7'b0000000, \
  7'b0000000 \
}

`define INIT_5x5_STATIC_BEEHIVE { \
  7'b0000000, \
  7'b0000000, \
  7'b0011000, \
  7'b0100100, \
  7'b0011000, \
  7'b0000000, \
  7'b0000000 \
}

`define INIT_5x5_STATIC_LOAF { \
  7'b0000000, \
  7'b0011000, \
  7'b0100100, \
  7'b0010100, \
  7'b0001000, \
  7'b0000000, \
  7'b0000000 \
}

`define INIT_5x5_STATIC_BOAT { \
  7'b0000000, \
  7'b0110000, \
  7'b0101000, \
  7'b0010000, \
  7'b0000000, \
  7'b0000000, \
  7'b0000000 \
}

`define INIT_5x5_STATIC_TUB { \
  7'b0000000, \
  7'b0000000, \
  7'b0001000, \
  7'b0010100, \
  7'b0001000, \
  7'b0000000, \
  7'b0000000 \
}

`define INIT_5x5_ALTERNATING { \
  7'b0000000, \
  7'b0101010, \
  7'b0010100, \
  7'b0101010, \
  7'b0010100, \
  7'b0101010, \
  7'b0000000 \
}

`define INIT_5x5_DBG1 { \
  7'b0000000, \
  7'b0001010, \
  7'b0000010, \
  7'b0010010, \
  7'b0000000, \
  7'b0000010, \
  7'b0000000 \
}

`define INIT_5x5_DBG2 { \
  7'b0000000, \
  7'b0010000, \
  7'b0000000, \
  7'b0100010, \
  7'b0000000, \
  7'b0001000, \
  7'b0000000 \
}


`define INIT_8x8_ALTERNATING { \
  10'b1010101010, \
  10'b0101010101, \
  10'b1010101010, \
  10'b0101010101, \
  10'b1010101010, \
  10'b0101010101, \
  10'b1010101010, \
  10'b0101010101, \
  10'b1010101010, \
  10'b0101010101 \
}

`define INIT_8x8_GLIDER { \
  10'b0000000000, \
  10'b0001000000, \
  10'b0000100000, \
  10'b0011100000, \
  10'b0000000000, \
  10'b0000000000, \
  10'b0000000000, \
  10'b0000000000, \
  10'b0000000000, \
  10'b0000000000 \
}


`define INIT_8x8_DIAGONAL { \
  10'b1000000000, \
  10'b0100000000, \
  10'b0010000000, \
  10'b0001000000, \
  10'b0000100000, \
  10'b0000010000, \
  10'b0000001000, \
  10'b0000000100, \
  10'b0000000010, \
  10'b0000000001 \
}


`define INIT_8x8_DOTS { \
  10'b0000000000, \
  10'b0100000000, \
  10'b0110000000, \
  10'b0111000000, \
  10'b0111100000, \
  10'b0111110000, \
  10'b0111111000, \
  10'b0111111100, \
  10'b0111111110, \
  10'b0000000000 \
}

`define INIT_8x8_FADING_BLINKERS { \
  10'b0000000000, \
  10'b0001110000, \
  10'b0000000000, \
  10'b0000000000, \
  10'b0001110000, \
  10'b0000000000, \
  10'b0000000000, \
  10'b0001110000, \
  10'b0000000000, \
  10'b0000000000 \
}

`define INIT_13x13_PULSAR { \
  17'b00000000000000000, \
  17'b00000000000000000, \
  17'b00001110001110000, \
  17'b00000000000000000, \
  17'b00100001010000100, \
  17'b00100001010000100, \
  17'b00100001010000100, \
  17'b00001110001110000, \
  17'b00000000000000000, \
  17'b00001110001110000, \
  17'b00100001010000100, \
  17'b00100001010000100, \
  17'b00100001010000100, \
  17'b00000000000000000, \
  17'b00001110001110000, \
  17'b00000000000000000, \
  17'b00000000000000000 \
}

`endif // INITIAL_CONDITIONS